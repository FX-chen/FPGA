module uart_rx(
    input sys_clk,
    input sys_rst_n,
    input uart_rxd,

    output reg uart_done,
    output reg [7:0] uart_data


);






endmodule